parameter RX_CFG = 14;
`define USE_WF
