parameter RX_CFG = 4;
`define USE_WF
