/*
--------------------------------------------------------------------------------
This library is free software; you can redistribute it and/or
modify it under the terms of the GNU Library General Public
License as published by the Free Software Foundation; either
version 2 of the License, or (at your option) any later version.
This library is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
Library General Public License for more details.
You should have received a copy of the GNU Library General Public
License along with this library; if not, write to the
Free Software Foundation, Inc., 51 Franklin St, Fifth Floor,
Boston, MA  02110-1301, USA.
--------------------------------------------------------------------------------
*/

// Copyright (c) 2008 Alex Shovkoplyas, VE3NEA
// Copyright (c) 2013 Phil Harman, VK6APH
// Copyright (c) 2014 John Seamons, ZL/KF6VO


// fixme: I can't remember the difference between cic_prune.v & cic_prune_var.v
// something about pre-shifting the input data?

//
// used in conjunction with .vh files generated by cic_gen.c
//
// implements 10-bit fixed (0-1024) and 5/10-bit 2**n variable decimation (R)
//
// NB: when variable decimation is specified by .DECIMATION(<0) then .GROWTH() must
// specify for the largest expected decimation.
//
// Fixed differential delay (D) = 1
//

module cic_prune (
	input wire clock,
	input wire reset,
	input wire [MD-1:0] decimation,
	input wire in_strobe,
	output reg out_strobe,
	input wire signed [IN_WIDTH-1:0] in_data,
	output reg signed [OUT_WIDTH-1:0] out_data
	);

	// design parameters
	parameter INCLUDE = "required";
	parameter DECIMATION = "required";  
	parameter GROWTH = "required";
	parameter IN_WIDTH = "required";
	parameter OUT_WIDTH = "required";
	
	localparam ACC_WIDTH = IN_WIDTH + GROWTH;

localparam MD = 13;		// max decim = 4096, assumes excess counter bits get optimized away

reg [MD-1:0] sample_no;
initial sample_no = {MD{1'b0}};
wire [MD-1:0] decim;

generate
	if (DECIMATION < 0) begin assign decim = decimation; end	// variable
	if (DECIMATION > 0) begin assign decim = DECIMATION; end	// fixed
endgenerate

always @(posedge clock)
  if (in_strobe)
    begin
    if (sample_no == (decim-1))
      begin
      sample_no <= 0;
      out_strobe <= 1;
      end
    else
      begin
      sample_no <= sample_no + 1'b1;
      out_strobe <= 0;
      end
    end
  else
    out_strobe <= 0;

wire signed [IN_WIDTH-1:0] in = in_data;
wire signed [OUT_WIDTH-1:0] out;

generate
	if (INCLUDE == "cic_rx1.vh") begin : rx1 `include "cic_rx1.vh" end
	if (INCLUDE == "cic_rx2.vh") begin : rx2 `include "cic_rx2.vh" end
	if (INCLUDE == "cic_wf1.vh") begin : wf1 `include "cic_wf1.vh" end
	if (INCLUDE == "cic_wf2.vh") begin : wf2 `include "cic_wf2.vh" end
endgenerate

generate
	if (DECIMATION < 0)
	begin
		always @(posedge clock)
			if (out_strobe)
				if (decim == 1)
					out_data <= in[IN_WIDTH-1 -:OUT_WIDTH];
				else
					out_data <= out;
	end
endgenerate

generate
	if (DECIMATION > 0)
	begin
		always @(posedge clock)
			if (out_strobe) out_data <= out;
	end
endgenerate

endmodule
