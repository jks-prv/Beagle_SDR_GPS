`ifndef _KIWI_VH_
`define _KIWI_VH_

// kiwi.inline.vh is appended by the e_cpu assembler to the generated file kiwi.gen.vh
// to make the new localparam scheme work

`endif
