localparam RX_CFG = 1;
`define USE_WF
