parameter RX_CFG = 4;
